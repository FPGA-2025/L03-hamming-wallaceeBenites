module calcula_hamming (
  input [10:0] entrada,
  output [14:0] saida
);

// implemente o seu código aqui

endmodule
